module W1_ROM (
    input  [2:0] addr,       // 0-31
    output reg signed [15:0] w1,
    output reg signed [15:0] w2,
    output reg signed [15:0] w3,
    output reg signed [15:0] w4
);

always @(*) begin

    // ---------------------- W1 ----------------------
    case (addr)
        0:  w1 = 28366;
        1:  w1 = 1235;
        2:  w1 = 32767;
        3:  w1 = 28311;
        4:  w1 = 27866;
        5:  w1 = -21901;
        6:  w1 = 11592;
        7:  w1 = -11250;
        default: w1 = 16'd0;
    endcase

    // ---------------------- W2 ----------------------
    case (addr)
        0:  w2 = -32768;
        1:  w2 = 7519;
        2:  w2 = 20296;
        3:  w2 = 11812;
        4:  w2 = 7880;
        5:  w2 = 11221;
        6:  w2 = 19840;
        7:  w2 = 9513;
        default: w2 = 16'd0;
    endcase

    // ---------------------- W3 ----------------------
    case (addr)
        0:  w3 = 20720;
        1:  w3 = -1834;
        2:  w3 = 19967;
        3:  w3 = -31414;
        4:  w3 = -32768;
        5:  w3 = -646;
        6:  w3 = 23343;
        7:  w3 = -16111;
        default: w3 = 16'd0;
    endcase

    // ---------------------- W4 ----------------------
    case (addr)
        0:  w4 = 32767;
        1:  w4 = -31614;
        2:  w4 = -32768;
        3:  w4 = 16909;
        4:  w4 = 30360;
        5:  w4 = 32767;
        6:  w4 = -5276;
        7:  w4 = 14196;
        default: w4 = 16'd0;
    endcase

end

endmodule
